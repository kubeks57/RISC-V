//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Sat Aug 10 20:24:59 2024
// Version: 2024.1 2024.1.0.3
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// M2_INTERFACE
module M2_INTERFACE(
    // Inputs
    ACLK,
    APB_TARGET_PADDR,
    APB_TARGET_PENABLE,
    APB_TARGET_PSEL,
    APB_TARGET_PWDATA,
    APB_TARGET_PWRITE,
    ARESETN,
    AXI4_INITIATOR_SLAVE0_ARREADY,
    AXI4_INITIATOR_SLAVE0_AWREADY,
    AXI4_INITIATOR_SLAVE0_BID,
    AXI4_INITIATOR_SLAVE0_BRESP,
    AXI4_INITIATOR_SLAVE0_BUSER,
    AXI4_INITIATOR_SLAVE0_BVALID,
    AXI4_INITIATOR_SLAVE0_RDATA,
    AXI4_INITIATOR_SLAVE0_RID,
    AXI4_INITIATOR_SLAVE0_RLAST,
    AXI4_INITIATOR_SLAVE0_RRESP,
    AXI4_INITIATOR_SLAVE0_RUSER,
    AXI4_INITIATOR_SLAVE0_RVALID,
    AXI4_INITIATOR_SLAVE0_WREADY,
    AXI_TARGET_MASTER0_ARADDR,
    AXI_TARGET_MASTER0_ARBURST,
    AXI_TARGET_MASTER0_ARCACHE,
    AXI_TARGET_MASTER0_ARID,
    AXI_TARGET_MASTER0_ARLEN,
    AXI_TARGET_MASTER0_ARLOCK,
    AXI_TARGET_MASTER0_ARPROT,
    AXI_TARGET_MASTER0_ARQOS,
    AXI_TARGET_MASTER0_ARREGION,
    AXI_TARGET_MASTER0_ARSIZE,
    AXI_TARGET_MASTER0_ARUSER,
    AXI_TARGET_MASTER0_ARVALID,
    AXI_TARGET_MASTER0_AWADDR,
    AXI_TARGET_MASTER0_AWBURST,
    AXI_TARGET_MASTER0_AWCACHE,
    AXI_TARGET_MASTER0_AWID,
    AXI_TARGET_MASTER0_AWLEN,
    AXI_TARGET_MASTER0_AWLOCK,
    AXI_TARGET_MASTER0_AWPROT,
    AXI_TARGET_MASTER0_AWQOS,
    AXI_TARGET_MASTER0_AWREGION,
    AXI_TARGET_MASTER0_AWSIZE,
    AXI_TARGET_MASTER0_AWUSER,
    AXI_TARGET_MASTER0_AWVALID,
    AXI_TARGET_MASTER0_BREADY,
    AXI_TARGET_MASTER0_RREADY,
    AXI_TARGET_MASTER0_WDATA,
    AXI_TARGET_MASTER0_WLAST,
    AXI_TARGET_MASTER0_WSTRB,
    AXI_TARGET_MASTER0_WUSER,
    AXI_TARGET_MASTER0_WVALID,
    CLKS_FROM_TXPLL_TO_PCIE_0_PCIE_0_TX_BIT_CLK,
    CLKS_FROM_TXPLL_TO_PCIE_0_PCIE_0_TX_PLL_LOCK,
    CLKS_FROM_TXPLL_TO_PCIE_0_PCIE_0_TX_PLL_REF_CLK,
    PCIESS_LANE_RXD0_N,
    PCIESS_LANE_RXD0_P,
    PCIE_0_TL_CLK_125MHz,
    PCIE_INIT_DONE,
    PCIE_REF_CLK,
    PCLK,
    PRESETN,
    // Outputs
    APB_TARGET_PRDATA,
    APB_TARGET_PREADY,
    APB_TARGET_PSLVERR,
    AXI4_INITIATOR_SLAVE0_ARADDR,
    AXI4_INITIATOR_SLAVE0_ARBURST,
    AXI4_INITIATOR_SLAVE0_ARCACHE,
    AXI4_INITIATOR_SLAVE0_ARID,
    AXI4_INITIATOR_SLAVE0_ARLEN,
    AXI4_INITIATOR_SLAVE0_ARLOCK,
    AXI4_INITIATOR_SLAVE0_ARPROT,
    AXI4_INITIATOR_SLAVE0_ARQOS,
    AXI4_INITIATOR_SLAVE0_ARREGION,
    AXI4_INITIATOR_SLAVE0_ARSIZE,
    AXI4_INITIATOR_SLAVE0_ARUSER,
    AXI4_INITIATOR_SLAVE0_ARVALID,
    AXI4_INITIATOR_SLAVE0_AWADDR,
    AXI4_INITIATOR_SLAVE0_AWBURST,
    AXI4_INITIATOR_SLAVE0_AWCACHE,
    AXI4_INITIATOR_SLAVE0_AWID,
    AXI4_INITIATOR_SLAVE0_AWLEN,
    AXI4_INITIATOR_SLAVE0_AWLOCK,
    AXI4_INITIATOR_SLAVE0_AWPROT,
    AXI4_INITIATOR_SLAVE0_AWQOS,
    AXI4_INITIATOR_SLAVE0_AWREGION,
    AXI4_INITIATOR_SLAVE0_AWSIZE,
    AXI4_INITIATOR_SLAVE0_AWUSER,
    AXI4_INITIATOR_SLAVE0_AWVALID,
    AXI4_INITIATOR_SLAVE0_BREADY,
    AXI4_INITIATOR_SLAVE0_RREADY,
    AXI4_INITIATOR_SLAVE0_WDATA,
    AXI4_INITIATOR_SLAVE0_WLAST,
    AXI4_INITIATOR_SLAVE0_WSTRB,
    AXI4_INITIATOR_SLAVE0_WUSER,
    AXI4_INITIATOR_SLAVE0_WVALID,
    AXI_TARGET_MASTER0_ARREADY,
    AXI_TARGET_MASTER0_AWREADY,
    AXI_TARGET_MASTER0_BID,
    AXI_TARGET_MASTER0_BRESP,
    AXI_TARGET_MASTER0_BUSER,
    AXI_TARGET_MASTER0_BVALID,
    AXI_TARGET_MASTER0_RDATA,
    AXI_TARGET_MASTER0_RID,
    AXI_TARGET_MASTER0_RLAST,
    AXI_TARGET_MASTER0_RRESP,
    AXI_TARGET_MASTER0_RUSER,
    AXI_TARGET_MASTER0_RVALID,
    AXI_TARGET_MASTER0_WREADY,
    M2_PERST0n,
    PCIESS_LANE_TXD0_N,
    PCIESS_LANE_TXD0_P,
    PCIE_INTERRUPT
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input         ACLK;
input  [25:0] APB_TARGET_PADDR;
input         APB_TARGET_PENABLE;
input         APB_TARGET_PSEL;
input  [31:0] APB_TARGET_PWDATA;
input         APB_TARGET_PWRITE;
input         ARESETN;
input         AXI4_INITIATOR_SLAVE0_ARREADY;
input         AXI4_INITIATOR_SLAVE0_AWREADY;
input  [4:0]  AXI4_INITIATOR_SLAVE0_BID;
input  [1:0]  AXI4_INITIATOR_SLAVE0_BRESP;
input  [0:0]  AXI4_INITIATOR_SLAVE0_BUSER;
input         AXI4_INITIATOR_SLAVE0_BVALID;
input  [63:0] AXI4_INITIATOR_SLAVE0_RDATA;
input  [4:0]  AXI4_INITIATOR_SLAVE0_RID;
input         AXI4_INITIATOR_SLAVE0_RLAST;
input  [1:0]  AXI4_INITIATOR_SLAVE0_RRESP;
input  [0:0]  AXI4_INITIATOR_SLAVE0_RUSER;
input         AXI4_INITIATOR_SLAVE0_RVALID;
input         AXI4_INITIATOR_SLAVE0_WREADY;
input  [37:0] AXI_TARGET_MASTER0_ARADDR;
input  [1:0]  AXI_TARGET_MASTER0_ARBURST;
input  [3:0]  AXI_TARGET_MASTER0_ARCACHE;
input  [7:0]  AXI_TARGET_MASTER0_ARID;
input  [7:0]  AXI_TARGET_MASTER0_ARLEN;
input  [1:0]  AXI_TARGET_MASTER0_ARLOCK;
input  [2:0]  AXI_TARGET_MASTER0_ARPROT;
input  [3:0]  AXI_TARGET_MASTER0_ARQOS;
input  [3:0]  AXI_TARGET_MASTER0_ARREGION;
input  [2:0]  AXI_TARGET_MASTER0_ARSIZE;
input  [0:0]  AXI_TARGET_MASTER0_ARUSER;
input         AXI_TARGET_MASTER0_ARVALID;
input  [37:0] AXI_TARGET_MASTER0_AWADDR;
input  [1:0]  AXI_TARGET_MASTER0_AWBURST;
input  [3:0]  AXI_TARGET_MASTER0_AWCACHE;
input  [7:0]  AXI_TARGET_MASTER0_AWID;
input  [7:0]  AXI_TARGET_MASTER0_AWLEN;
input  [1:0]  AXI_TARGET_MASTER0_AWLOCK;
input  [2:0]  AXI_TARGET_MASTER0_AWPROT;
input  [3:0]  AXI_TARGET_MASTER0_AWQOS;
input  [3:0]  AXI_TARGET_MASTER0_AWREGION;
input  [2:0]  AXI_TARGET_MASTER0_AWSIZE;
input  [0:0]  AXI_TARGET_MASTER0_AWUSER;
input         AXI_TARGET_MASTER0_AWVALID;
input         AXI_TARGET_MASTER0_BREADY;
input         AXI_TARGET_MASTER0_RREADY;
input  [63:0] AXI_TARGET_MASTER0_WDATA;
input         AXI_TARGET_MASTER0_WLAST;
input  [7:0]  AXI_TARGET_MASTER0_WSTRB;
input  [0:0]  AXI_TARGET_MASTER0_WUSER;
input         AXI_TARGET_MASTER0_WVALID;
input         CLKS_FROM_TXPLL_TO_PCIE_0_PCIE_0_TX_BIT_CLK;
input         CLKS_FROM_TXPLL_TO_PCIE_0_PCIE_0_TX_PLL_LOCK;
input         CLKS_FROM_TXPLL_TO_PCIE_0_PCIE_0_TX_PLL_REF_CLK;
input         PCIESS_LANE_RXD0_N;
input         PCIESS_LANE_RXD0_P;
input         PCIE_0_TL_CLK_125MHz;
input         PCIE_INIT_DONE;
input         PCIE_REF_CLK;
input         PCLK;
input         PRESETN;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [31:0] APB_TARGET_PRDATA;
output        APB_TARGET_PREADY;
output        APB_TARGET_PSLVERR;
output [37:0] AXI4_INITIATOR_SLAVE0_ARADDR;
output [1:0]  AXI4_INITIATOR_SLAVE0_ARBURST;
output [3:0]  AXI4_INITIATOR_SLAVE0_ARCACHE;
output [4:0]  AXI4_INITIATOR_SLAVE0_ARID;
output [7:0]  AXI4_INITIATOR_SLAVE0_ARLEN;
output [1:0]  AXI4_INITIATOR_SLAVE0_ARLOCK;
output [2:0]  AXI4_INITIATOR_SLAVE0_ARPROT;
output [3:0]  AXI4_INITIATOR_SLAVE0_ARQOS;
output [3:0]  AXI4_INITIATOR_SLAVE0_ARREGION;
output [2:0]  AXI4_INITIATOR_SLAVE0_ARSIZE;
output [0:0]  AXI4_INITIATOR_SLAVE0_ARUSER;
output        AXI4_INITIATOR_SLAVE0_ARVALID;
output [37:0] AXI4_INITIATOR_SLAVE0_AWADDR;
output [1:0]  AXI4_INITIATOR_SLAVE0_AWBURST;
output [3:0]  AXI4_INITIATOR_SLAVE0_AWCACHE;
output [4:0]  AXI4_INITIATOR_SLAVE0_AWID;
output [7:0]  AXI4_INITIATOR_SLAVE0_AWLEN;
output [1:0]  AXI4_INITIATOR_SLAVE0_AWLOCK;
output [2:0]  AXI4_INITIATOR_SLAVE0_AWPROT;
output [3:0]  AXI4_INITIATOR_SLAVE0_AWQOS;
output [3:0]  AXI4_INITIATOR_SLAVE0_AWREGION;
output [2:0]  AXI4_INITIATOR_SLAVE0_AWSIZE;
output [0:0]  AXI4_INITIATOR_SLAVE0_AWUSER;
output        AXI4_INITIATOR_SLAVE0_AWVALID;
output        AXI4_INITIATOR_SLAVE0_BREADY;
output        AXI4_INITIATOR_SLAVE0_RREADY;
output [63:0] AXI4_INITIATOR_SLAVE0_WDATA;
output        AXI4_INITIATOR_SLAVE0_WLAST;
output [7:0]  AXI4_INITIATOR_SLAVE0_WSTRB;
output [0:0]  AXI4_INITIATOR_SLAVE0_WUSER;
output        AXI4_INITIATOR_SLAVE0_WVALID;
output        AXI_TARGET_MASTER0_ARREADY;
output        AXI_TARGET_MASTER0_AWREADY;
output [7:0]  AXI_TARGET_MASTER0_BID;
output [1:0]  AXI_TARGET_MASTER0_BRESP;
output [0:0]  AXI_TARGET_MASTER0_BUSER;
output        AXI_TARGET_MASTER0_BVALID;
output [63:0] AXI_TARGET_MASTER0_RDATA;
output [7:0]  AXI_TARGET_MASTER0_RID;
output        AXI_TARGET_MASTER0_RLAST;
output [1:0]  AXI_TARGET_MASTER0_RRESP;
output [0:0]  AXI_TARGET_MASTER0_RUSER;
output        AXI_TARGET_MASTER0_RVALID;
output        AXI_TARGET_MASTER0_WREADY;
output        M2_PERST0n;
output        PCIESS_LANE_TXD0_N;
output        PCIESS_LANE_TXD0_P;
output        PCIE_INTERRUPT;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire          ACLK;
wire   [25:0] APB_TARGET_PADDR;
wire          APB_TARGET_PENABLE;
wire   [31:0] APB_TARGET_PRDATA_net_0;
wire          APB_TARGET_PREADY_net_0;
wire          APB_TARGET_PSEL;
wire          APB_TARGET_PSLVERR_net_0;
wire   [31:0] APB_TARGET_PWDATA;
wire          APB_TARGET_PWRITE;
wire          ARESETN;
wire   [37:0] AXI4_INITIATOR_ARADDR;
wire   [1:0]  AXI4_INITIATOR_ARBURST;
wire   [3:0]  AXI4_INITIATOR_ARCACHE;
wire   [4:0]  AXI4_INITIATOR_ARID;
wire   [7:0]  AXI4_INITIATOR_ARLEN;
wire   [1:0]  AXI4_INITIATOR_ARLOCK;
wire   [2:0]  AXI4_INITIATOR_ARPROT;
wire   [3:0]  AXI4_INITIATOR_ARQOS;
wire          AXI4_INITIATOR_SLAVE0_ARREADY;
wire   [3:0]  AXI4_INITIATOR_ARREGION;
wire   [2:0]  AXI4_INITIATOR_ARSIZE;
wire   [0:0]  AXI4_INITIATOR_ARUSER;
wire          AXI4_INITIATOR_ARVALID;
wire   [37:0] AXI4_INITIATOR_AWADDR;
wire   [1:0]  AXI4_INITIATOR_AWBURST;
wire   [3:0]  AXI4_INITIATOR_AWCACHE;
wire   [4:0]  AXI4_INITIATOR_AWID;
wire   [7:0]  AXI4_INITIATOR_AWLEN;
wire   [1:0]  AXI4_INITIATOR_AWLOCK;
wire   [2:0]  AXI4_INITIATOR_AWPROT;
wire   [3:0]  AXI4_INITIATOR_AWQOS;
wire          AXI4_INITIATOR_SLAVE0_AWREADY;
wire   [3:0]  AXI4_INITIATOR_AWREGION;
wire   [2:0]  AXI4_INITIATOR_AWSIZE;
wire   [0:0]  AXI4_INITIATOR_AWUSER;
wire          AXI4_INITIATOR_AWVALID;
wire   [4:0]  AXI4_INITIATOR_SLAVE0_BID;
wire          AXI4_INITIATOR_BREADY;
wire   [1:0]  AXI4_INITIATOR_SLAVE0_BRESP;
wire   [0:0]  AXI4_INITIATOR_SLAVE0_BUSER;
wire          AXI4_INITIATOR_SLAVE0_BVALID;
wire   [63:0] AXI4_INITIATOR_SLAVE0_RDATA;
wire   [4:0]  AXI4_INITIATOR_SLAVE0_RID;
wire          AXI4_INITIATOR_SLAVE0_RLAST;
wire          AXI4_INITIATOR_RREADY;
wire   [1:0]  AXI4_INITIATOR_SLAVE0_RRESP;
wire   [0:0]  AXI4_INITIATOR_SLAVE0_RUSER;
wire          AXI4_INITIATOR_SLAVE0_RVALID;
wire   [63:0] AXI4_INITIATOR_WDATA;
wire          AXI4_INITIATOR_WLAST;
wire          AXI4_INITIATOR_SLAVE0_WREADY;
wire   [7:0]  AXI4_INITIATOR_WSTRB;
wire   [0:0]  AXI4_INITIATOR_WUSER;
wire          AXI4_INITIATOR_WVALID;
wire   [37:0] AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARADDR;
wire   [1:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARBURST;
wire   [3:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARID;
wire   [7:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARLEN;
wire          AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARREADY;
wire          AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARVALID;
wire   [37:0] AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWADDR;
wire   [1:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWBURST;
wire   [3:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWID;
wire   [7:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWLEN;
wire          AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWREADY;
wire          AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWVALID;
wire   [3:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_BID;
wire          AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_BREADY;
wire   [1:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_BRESP;
wire   [0:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_BUSER;
wire          AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_BVALID;
wire   [63:0] AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RDATA;
wire   [3:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RID;
wire          AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RLAST;
wire          AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RREADY;
wire   [1:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RRESP;
wire   [0:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RUSER;
wire          AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RVALID;
wire   [63:0] AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WDATA;
wire          AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WLAST;
wire          AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WREADY;
wire   [7:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WSTRB;
wire          AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WVALID;
wire   [37:0] AXI_TARGET_MASTER0_ARADDR;
wire   [1:0]  AXI_TARGET_MASTER0_ARBURST;
wire   [3:0]  AXI_TARGET_MASTER0_ARCACHE;
wire   [7:0]  AXI_TARGET_MASTER0_ARID;
wire   [7:0]  AXI_TARGET_MASTER0_ARLEN;
wire   [1:0]  AXI_TARGET_MASTER0_ARLOCK;
wire   [2:0]  AXI_TARGET_MASTER0_ARPROT;
wire   [3:0]  AXI_TARGET_MASTER0_ARQOS;
wire          AXI_TARGET_ARREADY;
wire   [3:0]  AXI_TARGET_MASTER0_ARREGION;
wire   [2:0]  AXI_TARGET_MASTER0_ARSIZE;
wire   [0:0]  AXI_TARGET_MASTER0_ARUSER;
wire          AXI_TARGET_MASTER0_ARVALID;
wire   [37:0] AXI_TARGET_MASTER0_AWADDR;
wire   [1:0]  AXI_TARGET_MASTER0_AWBURST;
wire   [3:0]  AXI_TARGET_MASTER0_AWCACHE;
wire   [7:0]  AXI_TARGET_MASTER0_AWID;
wire   [7:0]  AXI_TARGET_MASTER0_AWLEN;
wire   [1:0]  AXI_TARGET_MASTER0_AWLOCK;
wire   [2:0]  AXI_TARGET_MASTER0_AWPROT;
wire   [3:0]  AXI_TARGET_MASTER0_AWQOS;
wire          AXI_TARGET_AWREADY;
wire   [3:0]  AXI_TARGET_MASTER0_AWREGION;
wire   [2:0]  AXI_TARGET_MASTER0_AWSIZE;
wire   [0:0]  AXI_TARGET_MASTER0_AWUSER;
wire          AXI_TARGET_MASTER0_AWVALID;
wire   [7:0]  AXI_TARGET_BID;
wire          AXI_TARGET_MASTER0_BREADY;
wire   [1:0]  AXI_TARGET_BRESP;
wire   [0:0]  AXI_TARGET_BUSER;
wire          AXI_TARGET_BVALID;
wire   [63:0] AXI_TARGET_RDATA;
wire   [7:0]  AXI_TARGET_RID;
wire          AXI_TARGET_RLAST;
wire          AXI_TARGET_MASTER0_RREADY;
wire   [1:0]  AXI_TARGET_RRESP;
wire   [0:0]  AXI_TARGET_RUSER;
wire          AXI_TARGET_RVALID;
wire   [63:0] AXI_TARGET_MASTER0_WDATA;
wire          AXI_TARGET_MASTER0_WLAST;
wire          AXI_TARGET_WREADY;
wire   [7:0]  AXI_TARGET_MASTER0_WSTRB;
wire   [0:0]  AXI_TARGET_MASTER0_WUSER;
wire          AXI_TARGET_MASTER0_WVALID;
wire          CLKS_FROM_TXPLL_TO_PCIE_0_PCIE_0_TX_BIT_CLK;
wire          CLKS_FROM_TXPLL_TO_PCIE_0_PCIE_0_TX_PLL_LOCK;
wire          CLKS_FROM_TXPLL_TO_PCIE_0_PCIE_0_TX_PLL_REF_CLK;
wire   [1:0]  FIC1_INITIATOR_AXI4mslave0_ARBURST;
wire   [3:0]  FIC1_INITIATOR_AXI4mslave0_ARCACHE;
wire   [7:0]  FIC1_INITIATOR_AXI4mslave0_ARLEN;
wire   [1:0]  FIC1_INITIATOR_AXI4mslave0_ARLOCK;
wire   [2:0]  FIC1_INITIATOR_AXI4mslave0_ARPROT;
wire   [3:0]  FIC1_INITIATOR_AXI4mslave0_ARQOS;
wire          FIC1_INITIATOR_AXI4mslave0_ARREADY;
wire   [3:0]  FIC1_INITIATOR_AXI4mslave0_ARREGION;
wire   [0:0]  FIC1_INITIATOR_AXI4mslave0_ARUSER;
wire          FIC1_INITIATOR_AXI4mslave0_ARVALID;
wire   [1:0]  FIC1_INITIATOR_AXI4mslave0_AWBURST;
wire   [3:0]  FIC1_INITIATOR_AXI4mslave0_AWCACHE;
wire   [7:0]  FIC1_INITIATOR_AXI4mslave0_AWLEN;
wire   [1:0]  FIC1_INITIATOR_AXI4mslave0_AWLOCK;
wire   [2:0]  FIC1_INITIATOR_AXI4mslave0_AWPROT;
wire   [3:0]  FIC1_INITIATOR_AXI4mslave0_AWQOS;
wire          FIC1_INITIATOR_AXI4mslave0_AWREADY;
wire   [3:0]  FIC1_INITIATOR_AXI4mslave0_AWREGION;
wire   [0:0]  FIC1_INITIATOR_AXI4mslave0_AWUSER;
wire          FIC1_INITIATOR_AXI4mslave0_AWVALID;
wire          FIC1_INITIATOR_AXI4mslave0_BREADY;
wire   [1:0]  FIC1_INITIATOR_AXI4mslave0_BRESP;
wire          FIC1_INITIATOR_AXI4mslave0_BVALID;
wire   [63:0] FIC1_INITIATOR_AXI4mslave0_RDATA;
wire          FIC1_INITIATOR_AXI4mslave0_RLAST;
wire          FIC1_INITIATOR_AXI4mslave0_RREADY;
wire   [1:0]  FIC1_INITIATOR_AXI4mslave0_RRESP;
wire          FIC1_INITIATOR_AXI4mslave0_RVALID;
wire   [63:0] FIC1_INITIATOR_AXI4mslave0_WDATA;
wire          FIC1_INITIATOR_AXI4mslave0_WLAST;
wire          FIC1_INITIATOR_AXI4mslave0_WREADY;
wire   [7:0]  FIC1_INITIATOR_AXI4mslave0_WSTRB;
wire   [0:0]  FIC1_INITIATOR_AXI4mslave0_WUSER;
wire          FIC1_INITIATOR_AXI4mslave0_WVALID;
wire          M2_PERST0n_net_0;
wire          PCIE_0_TL_CLK_125MHz;
wire   [31:0] PCIE_AXI_0_MASTER_ARADDR;
wire   [1:0]  PCIE_AXI_0_MASTER_ARBURST;
wire   [3:0]  PCIE_AXI_0_MASTER_ARID;
wire   [7:0]  PCIE_AXI_0_MASTER_ARLEN;
wire          PCIE_AXI_0_MASTER_ARREADY;
wire   [1:0]  PCIE_AXI_0_MASTER_ARSIZE;
wire          PCIE_AXI_0_MASTER_ARVALID;
wire   [31:0] PCIE_AXI_0_MASTER_AWADDR;
wire   [1:0]  PCIE_AXI_0_MASTER_AWBURST;
wire   [3:0]  PCIE_AXI_0_MASTER_AWID;
wire   [7:0]  PCIE_AXI_0_MASTER_AWLEN;
wire          PCIE_AXI_0_MASTER_AWREADY;
wire   [1:0]  PCIE_AXI_0_MASTER_AWSIZE;
wire          PCIE_AXI_0_MASTER_AWVALID;
wire   [3:0]  PCIE_AXI_0_MASTER_BID;
wire          PCIE_AXI_0_MASTER_BREADY;
wire   [1:0]  PCIE_AXI_0_MASTER_BRESP;
wire          PCIE_AXI_0_MASTER_BVALID;
wire   [63:0] PCIE_AXI_0_MASTER_RDATA;
wire   [3:0]  PCIE_AXI_0_MASTER_RID;
wire          PCIE_AXI_0_MASTER_RLAST;
wire          PCIE_AXI_0_MASTER_RREADY;
wire   [1:0]  PCIE_AXI_0_MASTER_RRESP;
wire          PCIE_AXI_0_MASTER_RVALID;
wire   [63:0] PCIE_AXI_0_MASTER_WDATA;
wire          PCIE_AXI_0_MASTER_WLAST;
wire          PCIE_AXI_0_MASTER_WREADY;
wire   [7:0]  PCIE_AXI_0_MASTER_WSTRB;
wire          PCIE_AXI_0_MASTER_WVALID;
wire          PCIE_INIT_DONE;
wire          PCIE_INTERRUPT_net_0;
wire          PCIE_REF_CLK;
wire          PCIESS_LANE_RXD0_N;
wire          PCIESS_LANE_RXD0_P;
wire          PCIESS_LANE_TXD0_N_net_0;
wire          PCIESS_LANE_TXD0_P_net_0;
wire          PCLK;
wire          PRESETN;
wire          APB_TARGET_PREADY_net_1;
wire          APB_TARGET_PSLVERR_net_1;
wire          AXI4_INITIATOR_ARVALID_net_0;
wire          AXI4_INITIATOR_AWVALID_net_0;
wire          AXI4_INITIATOR_BREADY_net_0;
wire          AXI4_INITIATOR_RREADY_net_0;
wire          AXI4_INITIATOR_WLAST_net_0;
wire          AXI4_INITIATOR_WVALID_net_0;
wire          AXI_TARGET_ARREADY_net_0;
wire          AXI_TARGET_AWREADY_net_0;
wire          AXI_TARGET_BVALID_net_0;
wire          AXI_TARGET_RLAST_net_0;
wire          AXI_TARGET_RVALID_net_0;
wire          AXI_TARGET_WREADY_net_0;
wire          M2_PERST0n_net_1;
wire          PCIESS_LANE_TXD0_N_net_1;
wire          PCIESS_LANE_TXD0_P_net_1;
wire          PCIE_INTERRUPT_net_1;
wire   [31:0] APB_TARGET_PRDATA_net_1;
wire   [37:0] AXI4_INITIATOR_ARADDR_net_0;
wire   [1:0]  AXI4_INITIATOR_ARBURST_net_0;
wire   [3:0]  AXI4_INITIATOR_ARCACHE_net_0;
wire   [4:0]  AXI4_INITIATOR_ARID_net_0;
wire   [7:0]  AXI4_INITIATOR_ARLEN_net_0;
wire   [1:0]  AXI4_INITIATOR_ARLOCK_net_0;
wire   [2:0]  AXI4_INITIATOR_ARPROT_net_0;
wire   [3:0]  AXI4_INITIATOR_ARQOS_net_0;
wire   [3:0]  AXI4_INITIATOR_ARREGION_net_0;
wire   [2:0]  AXI4_INITIATOR_ARSIZE_net_0;
wire   [0:0]  AXI4_INITIATOR_ARUSER_net_0;
wire   [37:0] AXI4_INITIATOR_AWADDR_net_0;
wire   [1:0]  AXI4_INITIATOR_AWBURST_net_0;
wire   [3:0]  AXI4_INITIATOR_AWCACHE_net_0;
wire   [4:0]  AXI4_INITIATOR_AWID_net_0;
wire   [7:0]  AXI4_INITIATOR_AWLEN_net_0;
wire   [1:0]  AXI4_INITIATOR_AWLOCK_net_0;
wire   [2:0]  AXI4_INITIATOR_AWPROT_net_0;
wire   [3:0]  AXI4_INITIATOR_AWQOS_net_0;
wire   [3:0]  AXI4_INITIATOR_AWREGION_net_0;
wire   [2:0]  AXI4_INITIATOR_AWSIZE_net_0;
wire   [0:0]  AXI4_INITIATOR_AWUSER_net_0;
wire   [63:0] AXI4_INITIATOR_WDATA_net_0;
wire   [7:0]  AXI4_INITIATOR_WSTRB_net_0;
wire   [0:0]  AXI4_INITIATOR_WUSER_net_0;
wire   [7:0]  AXI_TARGET_BID_net_0;
wire   [1:0]  AXI_TARGET_BRESP_net_0;
wire   [0:0]  AXI_TARGET_BUSER_net_0;
wire   [63:0] AXI_TARGET_RDATA_net_0;
wire   [7:0]  AXI_TARGET_RID_net_0;
wire   [1:0]  AXI_TARGET_RRESP_net_0;
wire   [0:0]  AXI_TARGET_RUSER_net_0;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire   [7:0]  PCIE_0_INTERRUPT_const_net_0;
wire          GND_net;
wire   [1:0]  MASTER0_AWLOCK_const_net_0;
wire   [3:0]  MASTER0_AWCACHE_const_net_0;
wire   [2:0]  MASTER0_AWPROT_const_net_0;
wire   [3:0]  MASTER0_AWQOS_const_net_0;
wire   [3:0]  MASTER0_AWREGION_const_net_0;
wire   [1:0]  MASTER0_ARLOCK_const_net_0;
wire   [3:0]  MASTER0_ARCACHE_const_net_0;
wire   [2:0]  MASTER0_ARPROT_const_net_0;
wire   [3:0]  MASTER0_ARQOS_const_net_0;
wire   [3:0]  MASTER0_ARREGION_const_net_0;
//--------------------------------------------------------------------
// Bus Interface Nets Declarations - Unequal Pin Widths
//--------------------------------------------------------------------
wire   [1:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARSIZE;
wire   [2:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARSIZE_0;
wire   [1:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARSIZE_0_1to0;
wire   [2:2]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARSIZE_0_2to2;
wire   [1:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWSIZE;
wire   [2:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWSIZE_0;
wire   [1:0]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWSIZE_0_1to0;
wire   [2:2]  AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWSIZE_0_2to2;
wire   [37:0] FIC1_INITIATOR_AXI4mslave0_ARADDR;
wire   [31:0] FIC1_INITIATOR_AXI4mslave0_ARADDR_0;
wire   [31:0] FIC1_INITIATOR_AXI4mslave0_ARADDR_0_31to0;
wire   [8:0]  FIC1_INITIATOR_AXI4mslave0_ARID;
wire   [3:0]  FIC1_INITIATOR_AXI4mslave0_ARID_0;
wire   [3:0]  FIC1_INITIATOR_AXI4mslave0_ARID_0_3to0;
wire   [2:0]  FIC1_INITIATOR_AXI4mslave0_ARSIZE;
wire   [1:0]  FIC1_INITIATOR_AXI4mslave0_ARSIZE_0;
wire   [1:0]  FIC1_INITIATOR_AXI4mslave0_ARSIZE_0_1to0;
wire   [37:0] FIC1_INITIATOR_AXI4mslave0_AWADDR;
wire   [31:0] FIC1_INITIATOR_AXI4mslave0_AWADDR_0;
wire   [31:0] FIC1_INITIATOR_AXI4mslave0_AWADDR_0_31to0;
wire   [8:0]  FIC1_INITIATOR_AXI4mslave0_AWID;
wire   [3:0]  FIC1_INITIATOR_AXI4mslave0_AWID_0;
wire   [3:0]  FIC1_INITIATOR_AXI4mslave0_AWID_0_3to0;
wire   [2:0]  FIC1_INITIATOR_AXI4mslave0_AWSIZE;
wire   [1:0]  FIC1_INITIATOR_AXI4mslave0_AWSIZE_0;
wire   [1:0]  FIC1_INITIATOR_AXI4mslave0_AWSIZE_0_1to0;
wire   [3:0]  FIC1_INITIATOR_AXI4mslave0_BID;
wire   [8:0]  FIC1_INITIATOR_AXI4mslave0_BID_0;
wire   [3:0]  FIC1_INITIATOR_AXI4mslave0_BID_0_3to0;
wire   [8:4]  FIC1_INITIATOR_AXI4mslave0_BID_0_8to4;
wire   [3:0]  FIC1_INITIATOR_AXI4mslave0_RID;
wire   [8:0]  FIC1_INITIATOR_AXI4mslave0_RID_0;
wire   [3:0]  FIC1_INITIATOR_AXI4mslave0_RID_0_3to0;
wire   [8:4]  FIC1_INITIATOR_AXI4mslave0_RID_0_8to4;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign PCIE_0_INTERRUPT_const_net_0 = 8'h00;
assign GND_net                      = 1'b0;
assign MASTER0_AWLOCK_const_net_0   = 2'h0;
assign MASTER0_AWCACHE_const_net_0  = 4'h0;
assign MASTER0_AWPROT_const_net_0   = 3'h0;
assign MASTER0_AWQOS_const_net_0    = 4'h0;
assign MASTER0_AWREGION_const_net_0 = 4'h0;
assign MASTER0_ARLOCK_const_net_0   = 2'h0;
assign MASTER0_ARCACHE_const_net_0  = 4'h0;
assign MASTER0_ARPROT_const_net_0   = 3'h0;
assign MASTER0_ARQOS_const_net_0    = 4'h0;
assign MASTER0_ARREGION_const_net_0 = 4'h0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign APB_TARGET_PREADY_net_1             = APB_TARGET_PREADY_net_0;
assign APB_TARGET_PREADY                   = APB_TARGET_PREADY_net_1;
assign APB_TARGET_PSLVERR_net_1            = APB_TARGET_PSLVERR_net_0;
assign APB_TARGET_PSLVERR                  = APB_TARGET_PSLVERR_net_1;
assign AXI4_INITIATOR_ARVALID_net_0        = AXI4_INITIATOR_ARVALID;
assign AXI4_INITIATOR_SLAVE0_ARVALID       = AXI4_INITIATOR_ARVALID_net_0;
assign AXI4_INITIATOR_AWVALID_net_0        = AXI4_INITIATOR_AWVALID;
assign AXI4_INITIATOR_SLAVE0_AWVALID       = AXI4_INITIATOR_AWVALID_net_0;
assign AXI4_INITIATOR_BREADY_net_0         = AXI4_INITIATOR_BREADY;
assign AXI4_INITIATOR_SLAVE0_BREADY        = AXI4_INITIATOR_BREADY_net_0;
assign AXI4_INITIATOR_RREADY_net_0         = AXI4_INITIATOR_RREADY;
assign AXI4_INITIATOR_SLAVE0_RREADY        = AXI4_INITIATOR_RREADY_net_0;
assign AXI4_INITIATOR_WLAST_net_0          = AXI4_INITIATOR_WLAST;
assign AXI4_INITIATOR_SLAVE0_WLAST         = AXI4_INITIATOR_WLAST_net_0;
assign AXI4_INITIATOR_WVALID_net_0         = AXI4_INITIATOR_WVALID;
assign AXI4_INITIATOR_SLAVE0_WVALID        = AXI4_INITIATOR_WVALID_net_0;
assign AXI_TARGET_ARREADY_net_0            = AXI_TARGET_ARREADY;
assign AXI_TARGET_MASTER0_ARREADY          = AXI_TARGET_ARREADY_net_0;
assign AXI_TARGET_AWREADY_net_0            = AXI_TARGET_AWREADY;
assign AXI_TARGET_MASTER0_AWREADY          = AXI_TARGET_AWREADY_net_0;
assign AXI_TARGET_BVALID_net_0             = AXI_TARGET_BVALID;
assign AXI_TARGET_MASTER0_BVALID           = AXI_TARGET_BVALID_net_0;
assign AXI_TARGET_RLAST_net_0              = AXI_TARGET_RLAST;
assign AXI_TARGET_MASTER0_RLAST            = AXI_TARGET_RLAST_net_0;
assign AXI_TARGET_RVALID_net_0             = AXI_TARGET_RVALID;
assign AXI_TARGET_MASTER0_RVALID           = AXI_TARGET_RVALID_net_0;
assign AXI_TARGET_WREADY_net_0             = AXI_TARGET_WREADY;
assign AXI_TARGET_MASTER0_WREADY           = AXI_TARGET_WREADY_net_0;
assign M2_PERST0n_net_1                    = M2_PERST0n_net_0;
assign M2_PERST0n                          = M2_PERST0n_net_1;
assign PCIESS_LANE_TXD0_N_net_1            = PCIESS_LANE_TXD0_N_net_0;
assign PCIESS_LANE_TXD0_N                  = PCIESS_LANE_TXD0_N_net_1;
assign PCIESS_LANE_TXD0_P_net_1            = PCIESS_LANE_TXD0_P_net_0;
assign PCIESS_LANE_TXD0_P                  = PCIESS_LANE_TXD0_P_net_1;
assign PCIE_INTERRUPT_net_1                = PCIE_INTERRUPT_net_0;
assign PCIE_INTERRUPT                      = PCIE_INTERRUPT_net_1;
assign APB_TARGET_PRDATA_net_1             = APB_TARGET_PRDATA_net_0;
assign APB_TARGET_PRDATA[31:0]             = APB_TARGET_PRDATA_net_1;
assign AXI4_INITIATOR_ARADDR_net_0         = AXI4_INITIATOR_ARADDR;
assign AXI4_INITIATOR_SLAVE0_ARADDR[37:0]  = AXI4_INITIATOR_ARADDR_net_0;
assign AXI4_INITIATOR_ARBURST_net_0        = AXI4_INITIATOR_ARBURST;
assign AXI4_INITIATOR_SLAVE0_ARBURST[1:0]  = AXI4_INITIATOR_ARBURST_net_0;
assign AXI4_INITIATOR_ARCACHE_net_0        = AXI4_INITIATOR_ARCACHE;
assign AXI4_INITIATOR_SLAVE0_ARCACHE[3:0]  = AXI4_INITIATOR_ARCACHE_net_0;
assign AXI4_INITIATOR_ARID_net_0           = AXI4_INITIATOR_ARID;
assign AXI4_INITIATOR_SLAVE0_ARID[4:0]     = AXI4_INITIATOR_ARID_net_0;
assign AXI4_INITIATOR_ARLEN_net_0          = AXI4_INITIATOR_ARLEN;
assign AXI4_INITIATOR_SLAVE0_ARLEN[7:0]    = AXI4_INITIATOR_ARLEN_net_0;
assign AXI4_INITIATOR_ARLOCK_net_0         = AXI4_INITIATOR_ARLOCK;
assign AXI4_INITIATOR_SLAVE0_ARLOCK[1:0]   = AXI4_INITIATOR_ARLOCK_net_0;
assign AXI4_INITIATOR_ARPROT_net_0         = AXI4_INITIATOR_ARPROT;
assign AXI4_INITIATOR_SLAVE0_ARPROT[2:0]   = AXI4_INITIATOR_ARPROT_net_0;
assign AXI4_INITIATOR_ARQOS_net_0          = AXI4_INITIATOR_ARQOS;
assign AXI4_INITIATOR_SLAVE0_ARQOS[3:0]    = AXI4_INITIATOR_ARQOS_net_0;
assign AXI4_INITIATOR_ARREGION_net_0       = AXI4_INITIATOR_ARREGION;
assign AXI4_INITIATOR_SLAVE0_ARREGION[3:0] = AXI4_INITIATOR_ARREGION_net_0;
assign AXI4_INITIATOR_ARSIZE_net_0         = AXI4_INITIATOR_ARSIZE;
assign AXI4_INITIATOR_SLAVE0_ARSIZE[2:0]   = AXI4_INITIATOR_ARSIZE_net_0;
assign AXI4_INITIATOR_ARUSER_net_0[0]      = AXI4_INITIATOR_ARUSER[0];
assign AXI4_INITIATOR_SLAVE0_ARUSER[0:0]   = AXI4_INITIATOR_ARUSER_net_0[0];
assign AXI4_INITIATOR_AWADDR_net_0         = AXI4_INITIATOR_AWADDR;
assign AXI4_INITIATOR_SLAVE0_AWADDR[37:0]  = AXI4_INITIATOR_AWADDR_net_0;
assign AXI4_INITIATOR_AWBURST_net_0        = AXI4_INITIATOR_AWBURST;
assign AXI4_INITIATOR_SLAVE0_AWBURST[1:0]  = AXI4_INITIATOR_AWBURST_net_0;
assign AXI4_INITIATOR_AWCACHE_net_0        = AXI4_INITIATOR_AWCACHE;
assign AXI4_INITIATOR_SLAVE0_AWCACHE[3:0]  = AXI4_INITIATOR_AWCACHE_net_0;
assign AXI4_INITIATOR_AWID_net_0           = AXI4_INITIATOR_AWID;
assign AXI4_INITIATOR_SLAVE0_AWID[4:0]     = AXI4_INITIATOR_AWID_net_0;
assign AXI4_INITIATOR_AWLEN_net_0          = AXI4_INITIATOR_AWLEN;
assign AXI4_INITIATOR_SLAVE0_AWLEN[7:0]    = AXI4_INITIATOR_AWLEN_net_0;
assign AXI4_INITIATOR_AWLOCK_net_0         = AXI4_INITIATOR_AWLOCK;
assign AXI4_INITIATOR_SLAVE0_AWLOCK[1:0]   = AXI4_INITIATOR_AWLOCK_net_0;
assign AXI4_INITIATOR_AWPROT_net_0         = AXI4_INITIATOR_AWPROT;
assign AXI4_INITIATOR_SLAVE0_AWPROT[2:0]   = AXI4_INITIATOR_AWPROT_net_0;
assign AXI4_INITIATOR_AWQOS_net_0          = AXI4_INITIATOR_AWQOS;
assign AXI4_INITIATOR_SLAVE0_AWQOS[3:0]    = AXI4_INITIATOR_AWQOS_net_0;
assign AXI4_INITIATOR_AWREGION_net_0       = AXI4_INITIATOR_AWREGION;
assign AXI4_INITIATOR_SLAVE0_AWREGION[3:0] = AXI4_INITIATOR_AWREGION_net_0;
assign AXI4_INITIATOR_AWSIZE_net_0         = AXI4_INITIATOR_AWSIZE;
assign AXI4_INITIATOR_SLAVE0_AWSIZE[2:0]   = AXI4_INITIATOR_AWSIZE_net_0;
assign AXI4_INITIATOR_AWUSER_net_0[0]      = AXI4_INITIATOR_AWUSER[0];
assign AXI4_INITIATOR_SLAVE0_AWUSER[0:0]   = AXI4_INITIATOR_AWUSER_net_0[0];
assign AXI4_INITIATOR_WDATA_net_0          = AXI4_INITIATOR_WDATA;
assign AXI4_INITIATOR_SLAVE0_WDATA[63:0]   = AXI4_INITIATOR_WDATA_net_0;
assign AXI4_INITIATOR_WSTRB_net_0          = AXI4_INITIATOR_WSTRB;
assign AXI4_INITIATOR_SLAVE0_WSTRB[7:0]    = AXI4_INITIATOR_WSTRB_net_0;
assign AXI4_INITIATOR_WUSER_net_0[0]       = AXI4_INITIATOR_WUSER[0];
assign AXI4_INITIATOR_SLAVE0_WUSER[0:0]    = AXI4_INITIATOR_WUSER_net_0[0];
assign AXI_TARGET_BID_net_0                = AXI_TARGET_BID;
assign AXI_TARGET_MASTER0_BID[7:0]         = AXI_TARGET_BID_net_0;
assign AXI_TARGET_BRESP_net_0              = AXI_TARGET_BRESP;
assign AXI_TARGET_MASTER0_BRESP[1:0]       = AXI_TARGET_BRESP_net_0;
assign AXI_TARGET_BUSER_net_0[0]           = AXI_TARGET_BUSER[0];
assign AXI_TARGET_MASTER0_BUSER[0:0]       = AXI_TARGET_BUSER_net_0[0];
assign AXI_TARGET_RDATA_net_0              = AXI_TARGET_RDATA;
assign AXI_TARGET_MASTER0_RDATA[63:0]      = AXI_TARGET_RDATA_net_0;
assign AXI_TARGET_RID_net_0                = AXI_TARGET_RID;
assign AXI_TARGET_MASTER0_RID[7:0]         = AXI_TARGET_RID_net_0;
assign AXI_TARGET_RRESP_net_0              = AXI_TARGET_RRESP;
assign AXI_TARGET_MASTER0_RRESP[1:0]       = AXI_TARGET_RRESP_net_0;
assign AXI_TARGET_RUSER_net_0[0]           = AXI_TARGET_RUSER[0];
assign AXI_TARGET_MASTER0_RUSER[0:0]       = AXI_TARGET_RUSER_net_0[0];
//--------------------------------------------------------------------
// Bus Interface Nets Assignments - Unequal Pin Widths
//--------------------------------------------------------------------
assign AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARSIZE_0 = { AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARSIZE_0_2to2, AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARSIZE_0_1to0 };
assign AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARSIZE_0_1to0 = AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARSIZE[1:0];
assign AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARSIZE_0_2to2 = 1'b0;

assign AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWSIZE_0 = { AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWSIZE_0_2to2, AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWSIZE_0_1to0 };
assign AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWSIZE_0_1to0 = AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWSIZE[1:0];
assign AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWSIZE_0_2to2 = 1'b0;

assign FIC1_INITIATOR_AXI4mslave0_ARADDR_0 = { FIC1_INITIATOR_AXI4mslave0_ARADDR_0_31to0 };
assign FIC1_INITIATOR_AXI4mslave0_ARADDR_0_31to0 = FIC1_INITIATOR_AXI4mslave0_ARADDR[31:0];

assign FIC1_INITIATOR_AXI4mslave0_ARID_0 = { FIC1_INITIATOR_AXI4mslave0_ARID_0_3to0 };
assign FIC1_INITIATOR_AXI4mslave0_ARID_0_3to0 = FIC1_INITIATOR_AXI4mslave0_ARID[3:0];

assign FIC1_INITIATOR_AXI4mslave0_ARSIZE_0 = { FIC1_INITIATOR_AXI4mslave0_ARSIZE_0_1to0 };
assign FIC1_INITIATOR_AXI4mslave0_ARSIZE_0_1to0 = FIC1_INITIATOR_AXI4mslave0_ARSIZE[1:0];

assign FIC1_INITIATOR_AXI4mslave0_AWADDR_0 = { FIC1_INITIATOR_AXI4mslave0_AWADDR_0_31to0 };
assign FIC1_INITIATOR_AXI4mslave0_AWADDR_0_31to0 = FIC1_INITIATOR_AXI4mslave0_AWADDR[31:0];

assign FIC1_INITIATOR_AXI4mslave0_AWID_0 = { FIC1_INITIATOR_AXI4mslave0_AWID_0_3to0 };
assign FIC1_INITIATOR_AXI4mslave0_AWID_0_3to0 = FIC1_INITIATOR_AXI4mslave0_AWID[3:0];

assign FIC1_INITIATOR_AXI4mslave0_AWSIZE_0 = { FIC1_INITIATOR_AXI4mslave0_AWSIZE_0_1to0 };
assign FIC1_INITIATOR_AXI4mslave0_AWSIZE_0_1to0 = FIC1_INITIATOR_AXI4mslave0_AWSIZE[1:0];

assign FIC1_INITIATOR_AXI4mslave0_BID_0 = { FIC1_INITIATOR_AXI4mslave0_BID_0_8to4, FIC1_INITIATOR_AXI4mslave0_BID_0_3to0 };
assign FIC1_INITIATOR_AXI4mslave0_BID_0_3to0 = FIC1_INITIATOR_AXI4mslave0_BID[3:0];
assign FIC1_INITIATOR_AXI4mslave0_BID_0_8to4 = 5'h0;

assign FIC1_INITIATOR_AXI4mslave0_RID_0 = { FIC1_INITIATOR_AXI4mslave0_RID_0_8to4, FIC1_INITIATOR_AXI4mslave0_RID_0_3to0 };
assign FIC1_INITIATOR_AXI4mslave0_RID_0_3to0 = FIC1_INITIATOR_AXI4mslave0_RID[3:0];
assign FIC1_INITIATOR_AXI4mslave0_RID_0_8to4 = 5'h0;

//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------AXI_ADDRESS_SHIM
AXI_ADDRESS_SHIM AXI_ADDRESS_SHIM_0(
        // Inputs
        .RESETN                ( ARESETN ),
        .INITIATOR_IN_ARREADY  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARREADY ),
        .INITIATOR_IN_AWREADY  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWREADY ),
        .INITIATOR_IN_BID      ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_BID ),
        .INITIATOR_IN_BRESP    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_BRESP ),
        .INITIATOR_IN_BVALID   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_BVALID ),
        .INITIATOR_IN_RDATA    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RDATA ),
        .INITIATOR_IN_RID      ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RID ),
        .INITIATOR_IN_RLAST    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RLAST ),
        .INITIATOR_IN_RRESP    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RRESP ),
        .INITIATOR_IN_RVALID   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RVALID ),
        .INITIATOR_IN_WREADY   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WREADY ),
        .TARGET_IN_ARADDR      ( PCIE_AXI_0_MASTER_ARADDR ),
        .TARGET_IN_ARBURST     ( PCIE_AXI_0_MASTER_ARBURST ),
        .TARGET_IN_ARID        ( PCIE_AXI_0_MASTER_ARID ),
        .TARGET_IN_ARLEN       ( PCIE_AXI_0_MASTER_ARLEN ),
        .TARGET_IN_ARSIZE      ( PCIE_AXI_0_MASTER_ARSIZE ),
        .TARGET_IN_ARVALID     ( PCIE_AXI_0_MASTER_ARVALID ),
        .TARGET_IN_AWADDR      ( PCIE_AXI_0_MASTER_AWADDR ),
        .TARGET_IN_AWBURST     ( PCIE_AXI_0_MASTER_AWBURST ),
        .TARGET_IN_AWID        ( PCIE_AXI_0_MASTER_AWID ),
        .TARGET_IN_AWLEN       ( PCIE_AXI_0_MASTER_AWLEN ),
        .TARGET_IN_AWSIZE      ( PCIE_AXI_0_MASTER_AWSIZE ),
        .TARGET_IN_AWVALID     ( PCIE_AXI_0_MASTER_AWVALID ),
        .TARGET_IN_BREADY      ( PCIE_AXI_0_MASTER_BREADY ),
        .TARGET_IN_RREADY      ( PCIE_AXI_0_MASTER_RREADY ),
        .TARGET_IN_WDATA       ( PCIE_AXI_0_MASTER_WDATA ),
        .TARGET_IN_WLAST       ( PCIE_AXI_0_MASTER_WLAST ),
        .TARGET_IN_WSTRB       ( PCIE_AXI_0_MASTER_WSTRB ),
        .TARGET_IN_WVALID      ( PCIE_AXI_0_MASTER_WVALID ),
        // Outputs
        .INITIATOR_OUT_ARADDR  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARADDR ),
        .INITIATOR_OUT_ARBURST ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARBURST ),
        .INITIATOR_OUT_ARID    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARID ),
        .INITIATOR_OUT_ARLEN   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARLEN ),
        .INITIATOR_OUT_ARSIZE  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARSIZE ),
        .INITIATOR_OUT_ARVALID ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARVALID ),
        .INITIATOR_OUT_AWADDR  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWADDR ),
        .INITIATOR_OUT_AWBURST ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWBURST ),
        .INITIATOR_OUT_AWID    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWID ),
        .INITIATOR_OUT_AWLEN   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWLEN ),
        .INITIATOR_OUT_AWSIZE  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWSIZE ),
        .INITIATOR_OUT_AWVALID ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWVALID ),
        .INITIATOR_OUT_BREADY  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_BREADY ),
        .INITIATOR_OUT_RREADY  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RREADY ),
        .INITIATOR_OUT_WDATA   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WDATA ),
        .INITIATOR_OUT_WLAST   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WLAST ),
        .INITIATOR_OUT_WSTRB   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WSTRB ),
        .INITIATOR_OUT_WVALID  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WVALID ),
        .TARGET_OUT_ARREADY    ( PCIE_AXI_0_MASTER_ARREADY ),
        .TARGET_OUT_AWREADY    ( PCIE_AXI_0_MASTER_AWREADY ),
        .TARGET_OUT_BID        ( PCIE_AXI_0_MASTER_BID ),
        .TARGET_OUT_BRESP      ( PCIE_AXI_0_MASTER_BRESP ),
        .TARGET_OUT_BVALID     ( PCIE_AXI_0_MASTER_BVALID ),
        .TARGET_OUT_RDATA      ( PCIE_AXI_0_MASTER_RDATA ),
        .TARGET_OUT_RID        ( PCIE_AXI_0_MASTER_RID ),
        .TARGET_OUT_RLAST      ( PCIE_AXI_0_MASTER_RLAST ),
        .TARGET_OUT_RRESP      ( PCIE_AXI_0_MASTER_RRESP ),
        .TARGET_OUT_RVALID     ( PCIE_AXI_0_MASTER_RVALID ),
        .TARGET_OUT_WREADY     ( PCIE_AXI_0_MASTER_WREADY ) 
        );

//--------FIC_1_INITIATOR
FIC_1_INITIATOR FIC1_INITIATOR(
        // Inputs
        .ACLK             ( ACLK ),
        .ARESETN          ( ARESETN ),
        .SLAVE0_AWREADY   ( FIC1_INITIATOR_AXI4mslave0_AWREADY ),
        .SLAVE0_WREADY    ( FIC1_INITIATOR_AXI4mslave0_WREADY ),
        .SLAVE0_BID       ( FIC1_INITIATOR_AXI4mslave0_BID_0 ),
        .SLAVE0_BRESP     ( FIC1_INITIATOR_AXI4mslave0_BRESP ),
        .SLAVE0_BVALID    ( FIC1_INITIATOR_AXI4mslave0_BVALID ),
        .SLAVE0_ARREADY   ( FIC1_INITIATOR_AXI4mslave0_ARREADY ),
        .SLAVE0_RID       ( FIC1_INITIATOR_AXI4mslave0_RID_0 ),
        .SLAVE0_RDATA     ( FIC1_INITIATOR_AXI4mslave0_RDATA ),
        .SLAVE0_RRESP     ( FIC1_INITIATOR_AXI4mslave0_RRESP ),
        .SLAVE0_RLAST     ( FIC1_INITIATOR_AXI4mslave0_RLAST ),
        .SLAVE0_RVALID    ( FIC1_INITIATOR_AXI4mslave0_RVALID ),
        .SLAVE0_BUSER     ( GND_net ), // tied to 1'b0 from definition
        .SLAVE0_RUSER     ( GND_net ), // tied to 1'b0 from definition
        .MASTER0_AWID     ( AXI_TARGET_MASTER0_AWID ),
        .MASTER0_AWADDR   ( AXI_TARGET_MASTER0_AWADDR ),
        .MASTER0_AWLEN    ( AXI_TARGET_MASTER0_AWLEN ),
        .MASTER0_AWSIZE   ( AXI_TARGET_MASTER0_AWSIZE ),
        .MASTER0_AWBURST  ( AXI_TARGET_MASTER0_AWBURST ),
        .MASTER0_AWLOCK   ( AXI_TARGET_MASTER0_AWLOCK ),
        .MASTER0_AWCACHE  ( AXI_TARGET_MASTER0_AWCACHE ),
        .MASTER0_AWPROT   ( AXI_TARGET_MASTER0_AWPROT ),
        .MASTER0_AWQOS    ( AXI_TARGET_MASTER0_AWQOS ),
        .MASTER0_AWREGION ( AXI_TARGET_MASTER0_AWREGION ),
        .MASTER0_AWVALID  ( AXI_TARGET_MASTER0_AWVALID ),
        .MASTER0_WDATA    ( AXI_TARGET_MASTER0_WDATA ),
        .MASTER0_WSTRB    ( AXI_TARGET_MASTER0_WSTRB ),
        .MASTER0_WLAST    ( AXI_TARGET_MASTER0_WLAST ),
        .MASTER0_WVALID   ( AXI_TARGET_MASTER0_WVALID ),
        .MASTER0_BREADY   ( AXI_TARGET_MASTER0_BREADY ),
        .MASTER0_ARID     ( AXI_TARGET_MASTER0_ARID ),
        .MASTER0_ARADDR   ( AXI_TARGET_MASTER0_ARADDR ),
        .MASTER0_ARLEN    ( AXI_TARGET_MASTER0_ARLEN ),
        .MASTER0_ARSIZE   ( AXI_TARGET_MASTER0_ARSIZE ),
        .MASTER0_ARBURST  ( AXI_TARGET_MASTER0_ARBURST ),
        .MASTER0_ARLOCK   ( AXI_TARGET_MASTER0_ARLOCK ),
        .MASTER0_ARCACHE  ( AXI_TARGET_MASTER0_ARCACHE ),
        .MASTER0_ARPROT   ( AXI_TARGET_MASTER0_ARPROT ),
        .MASTER0_ARQOS    ( AXI_TARGET_MASTER0_ARQOS ),
        .MASTER0_ARREGION ( AXI_TARGET_MASTER0_ARREGION ),
        .MASTER0_ARVALID  ( AXI_TARGET_MASTER0_ARVALID ),
        .MASTER0_RREADY   ( AXI_TARGET_MASTER0_RREADY ),
        .MASTER0_AWUSER   ( AXI_TARGET_MASTER0_AWUSER ),
        .MASTER0_WUSER    ( AXI_TARGET_MASTER0_WUSER ),
        .MASTER0_ARUSER   ( AXI_TARGET_MASTER0_ARUSER ),
        // Outputs
        .SLAVE0_AWID      ( FIC1_INITIATOR_AXI4mslave0_AWID ),
        .SLAVE0_AWADDR    ( FIC1_INITIATOR_AXI4mslave0_AWADDR ),
        .SLAVE0_AWLEN     ( FIC1_INITIATOR_AXI4mslave0_AWLEN ),
        .SLAVE0_AWSIZE    ( FIC1_INITIATOR_AXI4mslave0_AWSIZE ),
        .SLAVE0_AWBURST   ( FIC1_INITIATOR_AXI4mslave0_AWBURST ),
        .SLAVE0_AWLOCK    ( FIC1_INITIATOR_AXI4mslave0_AWLOCK ),
        .SLAVE0_AWCACHE   ( FIC1_INITIATOR_AXI4mslave0_AWCACHE ),
        .SLAVE0_AWPROT    ( FIC1_INITIATOR_AXI4mslave0_AWPROT ),
        .SLAVE0_AWQOS     ( FIC1_INITIATOR_AXI4mslave0_AWQOS ),
        .SLAVE0_AWREGION  ( FIC1_INITIATOR_AXI4mslave0_AWREGION ),
        .SLAVE0_AWVALID   ( FIC1_INITIATOR_AXI4mslave0_AWVALID ),
        .SLAVE0_WDATA     ( FIC1_INITIATOR_AXI4mslave0_WDATA ),
        .SLAVE0_WSTRB     ( FIC1_INITIATOR_AXI4mslave0_WSTRB ),
        .SLAVE0_WLAST     ( FIC1_INITIATOR_AXI4mslave0_WLAST ),
        .SLAVE0_WVALID    ( FIC1_INITIATOR_AXI4mslave0_WVALID ),
        .SLAVE0_BREADY    ( FIC1_INITIATOR_AXI4mslave0_BREADY ),
        .SLAVE0_ARID      ( FIC1_INITIATOR_AXI4mslave0_ARID ),
        .SLAVE0_ARADDR    ( FIC1_INITIATOR_AXI4mslave0_ARADDR ),
        .SLAVE0_ARLEN     ( FIC1_INITIATOR_AXI4mslave0_ARLEN ),
        .SLAVE0_ARSIZE    ( FIC1_INITIATOR_AXI4mslave0_ARSIZE ),
        .SLAVE0_ARBURST   ( FIC1_INITIATOR_AXI4mslave0_ARBURST ),
        .SLAVE0_ARLOCK    ( FIC1_INITIATOR_AXI4mslave0_ARLOCK ),
        .SLAVE0_ARCACHE   ( FIC1_INITIATOR_AXI4mslave0_ARCACHE ),
        .SLAVE0_ARPROT    ( FIC1_INITIATOR_AXI4mslave0_ARPROT ),
        .SLAVE0_ARQOS     ( FIC1_INITIATOR_AXI4mslave0_ARQOS ),
        .SLAVE0_ARREGION  ( FIC1_INITIATOR_AXI4mslave0_ARREGION ),
        .SLAVE0_ARVALID   ( FIC1_INITIATOR_AXI4mslave0_ARVALID ),
        .SLAVE0_RREADY    ( FIC1_INITIATOR_AXI4mslave0_RREADY ),
        .SLAVE0_AWUSER    ( FIC1_INITIATOR_AXI4mslave0_AWUSER ),
        .SLAVE0_WUSER     ( FIC1_INITIATOR_AXI4mslave0_WUSER ),
        .SLAVE0_ARUSER    ( FIC1_INITIATOR_AXI4mslave0_ARUSER ),
        .MASTER0_AWREADY  ( AXI_TARGET_AWREADY ),
        .MASTER0_WREADY   ( AXI_TARGET_WREADY ),
        .MASTER0_BID      ( AXI_TARGET_BID ),
        .MASTER0_BRESP    ( AXI_TARGET_BRESP ),
        .MASTER0_BVALID   ( AXI_TARGET_BVALID ),
        .MASTER0_ARREADY  ( AXI_TARGET_ARREADY ),
        .MASTER0_RID      ( AXI_TARGET_RID ),
        .MASTER0_RDATA    ( AXI_TARGET_RDATA ),
        .MASTER0_RRESP    ( AXI_TARGET_RRESP ),
        .MASTER0_RLAST    ( AXI_TARGET_RLAST ),
        .MASTER0_RVALID   ( AXI_TARGET_RVALID ),
        .MASTER0_BUSER    ( AXI_TARGET_BUSER ),
        .MASTER0_RUSER    ( AXI_TARGET_RUSER ) 
        );

//--------PF_PCIE_C0
PF_PCIE_C0 PCIE(
        // Inputs
        .INIT_DONE                  ( PCIE_INIT_DONE ),
        .APB_S_PRESET_N             ( PRESETN ),
        .APB_S_PCLK                 ( PCLK ),
        .PCIESS_AXI_0_S_ARBURST     ( FIC1_INITIATOR_AXI4mslave0_ARBURST ),
        .PCIESS_AXI_0_S_ARID        ( FIC1_INITIATOR_AXI4mslave0_ARID_0 ),
        .PCIESS_AXI_0_S_ARLEN       ( FIC1_INITIATOR_AXI4mslave0_ARLEN ),
        .PCIESS_AXI_0_S_ARSIZE      ( FIC1_INITIATOR_AXI4mslave0_ARSIZE_0 ),
        .PCIESS_AXI_0_S_ARVALID     ( FIC1_INITIATOR_AXI4mslave0_ARVALID ),
        .PCIESS_AXI_0_S_AWBURST     ( FIC1_INITIATOR_AXI4mslave0_AWBURST ),
        .PCIESS_AXI_0_S_AWID        ( FIC1_INITIATOR_AXI4mslave0_AWID_0 ),
        .PCIESS_AXI_0_S_AWLEN       ( FIC1_INITIATOR_AXI4mslave0_AWLEN ),
        .PCIESS_AXI_0_S_AWSIZE      ( FIC1_INITIATOR_AXI4mslave0_AWSIZE_0 ),
        .PCIESS_AXI_0_S_AWVALID     ( FIC1_INITIATOR_AXI4mslave0_AWVALID ),
        .PCIESS_AXI_0_S_BREADY      ( FIC1_INITIATOR_AXI4mslave0_BREADY ),
        .PCIESS_AXI_0_S_RREADY      ( FIC1_INITIATOR_AXI4mslave0_RREADY ),
        .PCIESS_AXI_0_S_WSTRB       ( FIC1_INITIATOR_AXI4mslave0_WSTRB ),
        .PCIESS_AXI_0_S_WLAST       ( FIC1_INITIATOR_AXI4mslave0_WLAST ),
        .PCIESS_AXI_0_S_WVALID      ( FIC1_INITIATOR_AXI4mslave0_WVALID ),
        .PCIESS_AXI_0_S_AWADDR      ( FIC1_INITIATOR_AXI4mslave0_AWADDR_0 ),
        .PCIESS_AXI_0_S_WDATA       ( FIC1_INITIATOR_AXI4mslave0_WDATA ),
        .PCIESS_AXI_0_S_ARADDR      ( FIC1_INITIATOR_AXI4mslave0_ARADDR_0 ),
        .PCIESS_AXI_0_M_ARREADY     ( PCIE_AXI_0_MASTER_ARREADY ),
        .PCIESS_AXI_0_M_AWREADY     ( PCIE_AXI_0_MASTER_AWREADY ),
        .PCIESS_AXI_0_M_BID         ( PCIE_AXI_0_MASTER_BID ),
        .PCIESS_AXI_0_M_BRESP       ( PCIE_AXI_0_MASTER_BRESP ),
        .PCIESS_AXI_0_M_BVALID      ( PCIE_AXI_0_MASTER_BVALID ),
        .PCIESS_AXI_0_M_RID         ( PCIE_AXI_0_MASTER_RID ),
        .PCIESS_AXI_0_M_RRESP       ( PCIE_AXI_0_MASTER_RRESP ),
        .PCIESS_AXI_0_M_RLAST       ( PCIE_AXI_0_MASTER_RLAST ),
        .PCIESS_AXI_0_M_RVALID      ( PCIE_AXI_0_MASTER_RVALID ),
        .PCIESS_AXI_0_M_WREADY      ( PCIE_AXI_0_MASTER_WREADY ),
        .PCIESS_AXI_0_M_RDATA       ( PCIE_AXI_0_MASTER_RDATA ),
        .APB_S_PSEL                 ( APB_TARGET_PSEL ),
        .APB_S_PENABLE              ( APB_TARGET_PENABLE ),
        .APB_S_PWRITE               ( APB_TARGET_PWRITE ),
        .APB_S_PADDR                ( APB_TARGET_PADDR ),
        .APB_S_PWDATA               ( APB_TARGET_PWDATA ),
        .PCIE_0_TX_PLL_LOCK         ( CLKS_FROM_TXPLL_TO_PCIE_0_PCIE_0_TX_PLL_LOCK ),
        .PCIE_0_TX_BIT_CLK          ( CLKS_FROM_TXPLL_TO_PCIE_0_PCIE_0_TX_BIT_CLK ),
        .PCIE_0_TX_PLL_REF_CLK      ( CLKS_FROM_TXPLL_TO_PCIE_0_PCIE_0_TX_PLL_REF_CLK ),
        .PCIESS_LANE_RXD0_P         ( PCIESS_LANE_RXD0_P ),
        .PCIESS_LANE_RXD0_N         ( PCIESS_LANE_RXD0_N ),
        .PCIESS_LANE0_CDR_REF_CLK_0 ( PCIE_REF_CLK ),
        .AXI_CLK                    ( ACLK ),
        .AXI_CLK_STABLE             ( ARESETN ),
        .PCIE_0_TL_CLK_125MHz       ( PCIE_0_TL_CLK_125MHz ),
        .PCIE_0_INTERRUPT           ( PCIE_0_INTERRUPT_const_net_0 ),
        .PCIE_0_M_RDERR             ( GND_net ),
        .PCIE_0_S_WDERR             ( GND_net ),
        // Outputs
        .PCIESS_AXI_0_S_ARREADY     ( FIC1_INITIATOR_AXI4mslave0_ARREADY ),
        .PCIESS_AXI_0_S_AWREADY     ( FIC1_INITIATOR_AXI4mslave0_AWREADY ),
        .PCIESS_AXI_0_S_BID         ( FIC1_INITIATOR_AXI4mslave0_BID ),
        .PCIESS_AXI_0_S_BRESP       ( FIC1_INITIATOR_AXI4mslave0_BRESP ),
        .PCIESS_AXI_0_S_BVALID      ( FIC1_INITIATOR_AXI4mslave0_BVALID ),
        .PCIESS_AXI_0_S_RID         ( FIC1_INITIATOR_AXI4mslave0_RID ),
        .PCIESS_AXI_0_S_RRESP       ( FIC1_INITIATOR_AXI4mslave0_RRESP ),
        .PCIESS_AXI_0_S_RLAST       ( FIC1_INITIATOR_AXI4mslave0_RLAST ),
        .PCIESS_AXI_0_S_RVALID      ( FIC1_INITIATOR_AXI4mslave0_RVALID ),
        .PCIESS_AXI_0_S_WREADY      ( FIC1_INITIATOR_AXI4mslave0_WREADY ),
        .PCIESS_AXI_0_S_RDATA       ( FIC1_INITIATOR_AXI4mslave0_RDATA ),
        .PCIESS_AXI_0_M_ARBURST     ( PCIE_AXI_0_MASTER_ARBURST ),
        .PCIESS_AXI_0_M_ARLEN       ( PCIE_AXI_0_MASTER_ARLEN ),
        .PCIESS_AXI_0_M_ARSIZE      ( PCIE_AXI_0_MASTER_ARSIZE ),
        .PCIESS_AXI_0_M_ARVALID     ( PCIE_AXI_0_MASTER_ARVALID ),
        .PCIESS_AXI_0_M_AWBURST     ( PCIE_AXI_0_MASTER_AWBURST ),
        .PCIESS_AXI_0_M_AWLEN       ( PCIE_AXI_0_MASTER_AWLEN ),
        .PCIESS_AXI_0_M_AWSIZE      ( PCIE_AXI_0_MASTER_AWSIZE ),
        .PCIESS_AXI_0_M_AWVALID     ( PCIE_AXI_0_MASTER_AWVALID ),
        .PCIESS_AXI_0_M_BREADY      ( PCIE_AXI_0_MASTER_BREADY ),
        .PCIESS_AXI_0_M_RREADY      ( PCIE_AXI_0_MASTER_RREADY ),
        .PCIESS_AXI_0_M_WSTRB       ( PCIE_AXI_0_MASTER_WSTRB ),
        .PCIESS_AXI_0_M_WLAST       ( PCIE_AXI_0_MASTER_WLAST ),
        .PCIESS_AXI_0_M_WVALID      ( PCIE_AXI_0_MASTER_WVALID ),
        .PCIESS_AXI_0_M_ARID        ( PCIE_AXI_0_MASTER_ARID ),
        .PCIESS_AXI_0_M_AWADDR      ( PCIE_AXI_0_MASTER_AWADDR ),
        .PCIESS_AXI_0_M_WDATA       ( PCIE_AXI_0_MASTER_WDATA ),
        .PCIESS_AXI_0_M_AWID        ( PCIE_AXI_0_MASTER_AWID ),
        .PCIESS_AXI_0_M_ARADDR      ( PCIE_AXI_0_MASTER_ARADDR ),
        .APB_S_PREADY               ( APB_TARGET_PREADY_net_0 ),
        .APB_S_PRDATA               ( APB_TARGET_PRDATA_net_0 ),
        .APB_S_PSLVERR              ( APB_TARGET_PSLVERR_net_0 ),
        .PCIESS_LANE_TXD0_P         ( PCIESS_LANE_TXD0_P_net_0 ),
        .PCIESS_LANE_TXD0_N         ( PCIESS_LANE_TXD0_N_net_0 ),
        .PCIE_0_LTSSM               (  ),
        .PCIE_0_INTERRUPT_OUT       ( PCIE_INTERRUPT_net_0 ),
        .PCIE_0_M_WDERR             (  ),
        .PCIE_0_S_RDERR             (  ),
        .PCIE_0_HOT_RST_EXIT        (  ),
        .PCIE_0_DLUP_EXIT           (  ),
        .PCIE_0_PERST_OUT_N         ( M2_PERST0n_net_0 ) 
        );

//--------PCIE_INITIATOR
PCIE_INITIATOR PCIE_INITIATOR_inst_0(
        // Inputs
        .ACLK             ( ACLK ),
        .ARESETN          ( ARESETN ),
        .SLAVE0_AWREADY   ( AXI4_INITIATOR_SLAVE0_AWREADY ),
        .SLAVE0_WREADY    ( AXI4_INITIATOR_SLAVE0_WREADY ),
        .SLAVE0_BID       ( AXI4_INITIATOR_SLAVE0_BID ),
        .SLAVE0_BRESP     ( AXI4_INITIATOR_SLAVE0_BRESP ),
        .SLAVE0_BVALID    ( AXI4_INITIATOR_SLAVE0_BVALID ),
        .SLAVE0_ARREADY   ( AXI4_INITIATOR_SLAVE0_ARREADY ),
        .SLAVE0_RID       ( AXI4_INITIATOR_SLAVE0_RID ),
        .SLAVE0_RDATA     ( AXI4_INITIATOR_SLAVE0_RDATA ),
        .SLAVE0_RRESP     ( AXI4_INITIATOR_SLAVE0_RRESP ),
        .SLAVE0_RLAST     ( AXI4_INITIATOR_SLAVE0_RLAST ),
        .SLAVE0_RVALID    ( AXI4_INITIATOR_SLAVE0_RVALID ),
        .SLAVE0_BUSER     ( AXI4_INITIATOR_SLAVE0_BUSER ),
        .SLAVE0_RUSER     ( AXI4_INITIATOR_SLAVE0_RUSER ),
        .MASTER0_AWID     ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWID ),
        .MASTER0_AWADDR   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWADDR ),
        .MASTER0_AWLEN    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWLEN ),
        .MASTER0_AWSIZE   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWSIZE_0 ),
        .MASTER0_AWBURST  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWBURST ),
        .MASTER0_AWLOCK   ( MASTER0_AWLOCK_const_net_0 ), // tied to 2'h0 from definition
        .MASTER0_AWCACHE  ( MASTER0_AWCACHE_const_net_0 ), // tied to 4'h0 from definition
        .MASTER0_AWPROT   ( MASTER0_AWPROT_const_net_0 ), // tied to 3'h0 from definition
        .MASTER0_AWQOS    ( MASTER0_AWQOS_const_net_0 ), // tied to 4'h0 from definition
        .MASTER0_AWREGION ( MASTER0_AWREGION_const_net_0 ), // tied to 4'h0 from definition
        .MASTER0_AWVALID  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWVALID ),
        .MASTER0_WDATA    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WDATA ),
        .MASTER0_WSTRB    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WSTRB ),
        .MASTER0_WLAST    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WLAST ),
        .MASTER0_WVALID   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WVALID ),
        .MASTER0_BREADY   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_BREADY ),
        .MASTER0_ARID     ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARID ),
        .MASTER0_ARADDR   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARADDR ),
        .MASTER0_ARLEN    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARLEN ),
        .MASTER0_ARSIZE   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARSIZE_0 ),
        .MASTER0_ARBURST  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARBURST ),
        .MASTER0_ARLOCK   ( MASTER0_ARLOCK_const_net_0 ), // tied to 2'h0 from definition
        .MASTER0_ARCACHE  ( MASTER0_ARCACHE_const_net_0 ), // tied to 4'h0 from definition
        .MASTER0_ARPROT   ( MASTER0_ARPROT_const_net_0 ), // tied to 3'h0 from definition
        .MASTER0_ARQOS    ( MASTER0_ARQOS_const_net_0 ), // tied to 4'h0 from definition
        .MASTER0_ARREGION ( MASTER0_ARREGION_const_net_0 ), // tied to 4'h0 from definition
        .MASTER0_ARVALID  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARVALID ),
        .MASTER0_RREADY   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RREADY ),
        .MASTER0_AWUSER   ( GND_net ), // tied to 1'b0 from definition
        .MASTER0_WUSER    ( GND_net ), // tied to 1'b0 from definition
        .MASTER0_ARUSER   ( GND_net ), // tied to 1'b0 from definition
        // Outputs
        .SLAVE0_AWID      ( AXI4_INITIATOR_AWID ),
        .SLAVE0_AWADDR    ( AXI4_INITIATOR_AWADDR ),
        .SLAVE0_AWLEN     ( AXI4_INITIATOR_AWLEN ),
        .SLAVE0_AWSIZE    ( AXI4_INITIATOR_AWSIZE ),
        .SLAVE0_AWBURST   ( AXI4_INITIATOR_AWBURST ),
        .SLAVE0_AWLOCK    ( AXI4_INITIATOR_AWLOCK ),
        .SLAVE0_AWCACHE   ( AXI4_INITIATOR_AWCACHE ),
        .SLAVE0_AWPROT    ( AXI4_INITIATOR_AWPROT ),
        .SLAVE0_AWQOS     ( AXI4_INITIATOR_AWQOS ),
        .SLAVE0_AWREGION  ( AXI4_INITIATOR_AWREGION ),
        .SLAVE0_AWVALID   ( AXI4_INITIATOR_AWVALID ),
        .SLAVE0_WDATA     ( AXI4_INITIATOR_WDATA ),
        .SLAVE0_WSTRB     ( AXI4_INITIATOR_WSTRB ),
        .SLAVE0_WLAST     ( AXI4_INITIATOR_WLAST ),
        .SLAVE0_WVALID    ( AXI4_INITIATOR_WVALID ),
        .SLAVE0_BREADY    ( AXI4_INITIATOR_BREADY ),
        .SLAVE0_ARID      ( AXI4_INITIATOR_ARID ),
        .SLAVE0_ARADDR    ( AXI4_INITIATOR_ARADDR ),
        .SLAVE0_ARLEN     ( AXI4_INITIATOR_ARLEN ),
        .SLAVE0_ARSIZE    ( AXI4_INITIATOR_ARSIZE ),
        .SLAVE0_ARBURST   ( AXI4_INITIATOR_ARBURST ),
        .SLAVE0_ARLOCK    ( AXI4_INITIATOR_ARLOCK ),
        .SLAVE0_ARCACHE   ( AXI4_INITIATOR_ARCACHE ),
        .SLAVE0_ARPROT    ( AXI4_INITIATOR_ARPROT ),
        .SLAVE0_ARQOS     ( AXI4_INITIATOR_ARQOS ),
        .SLAVE0_ARREGION  ( AXI4_INITIATOR_ARREGION ),
        .SLAVE0_ARVALID   ( AXI4_INITIATOR_ARVALID ),
        .SLAVE0_RREADY    ( AXI4_INITIATOR_RREADY ),
        .SLAVE0_AWUSER    ( AXI4_INITIATOR_AWUSER ),
        .SLAVE0_WUSER     ( AXI4_INITIATOR_WUSER ),
        .SLAVE0_ARUSER    ( AXI4_INITIATOR_ARUSER ),
        .MASTER0_AWREADY  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_AWREADY ),
        .MASTER0_WREADY   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_WREADY ),
        .MASTER0_BID      ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_BID ),
        .MASTER0_BRESP    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_BRESP ),
        .MASTER0_BVALID   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_BVALID ),
        .MASTER0_ARREADY  ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_ARREADY ),
        .MASTER0_RID      ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RID ),
        .MASTER0_RDATA    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RDATA ),
        .MASTER0_RRESP    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RRESP ),
        .MASTER0_RLAST    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RLAST ),
        .MASTER0_RVALID   ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RVALID ),
        .MASTER0_BUSER    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_BUSER ),
        .MASTER0_RUSER    ( AXI_ADDRESS_SHIM_0_AXI4_INITIATOR_RUSER ) 
        );


endmodule
